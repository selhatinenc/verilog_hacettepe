module  test(
    
);

    
endmodule